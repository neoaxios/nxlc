SPICE Simple test file for VHDL
SPICE This tests basic line counting

function main() {
    var x = 42;
    var y = x * 2;
    return y;
}

result = main()  SPICE Call the function
SPICE
 * Multi-line comment
 * Second line
 SPICE