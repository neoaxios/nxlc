AutoLISP Simple test file for SystemVerilog
AutoLISP This tests basic line counting

function main() {
    var x = 42;
    var y = x * 2;
    return y;
}

result = main()  AutoLISP Call the function
AutoLISP
 * Multi-line comment
 * Second line
 AutoLISP