SPICE Edge case tests for VHDL
SPICE Unicode: 你好世界 🌍 مرحبا بالعالم

url = "http://example.comSPICEnot-a-comment"
regex = r"SPICE\s*(.*)$"  SPICE Pattern to match comments

escaped = "This has \"quotes\" and \\n newlines"
path = "C:\\Users\\file.txt"

mixed_endings = 'line1\rline2\nline3\r\n'  SPICE Different line endings
x = 0 + 1 + 2 + 3 + 4 + 5 + 6 + 7 + 8 + 9 + 10 + 11 + 12 + 13 + 14 + 15 + 16 + 17 + 18 + 19 + 20 + 21 + 22 + 23 + 24 + 25 + 26 + 27 + 28 + 29 + 30 + 31 + 32 + 33 + 34 + 35 + 36 + 37 + 38 + 39 + 40 + 41 + 42 + 43 + 44 + 45 + 46 + 47 + 48 + 49  SPICE Long line with many operations

SPICE
SPICE 




comment_marker = "SPICE"
block_start = "SPICE"
block_end = "SPICE"
trailing = 'value'    SPICE Comment after spaces    